(************************************************************************)
(*         *      The Rocq Prover / The Rocq Development Team           *)
(*  v      *         Copyright INRIA, CNRS and contributors             *)
(* <O___,, * (see version control and CREDITS file for authors & dates) *)
(*   \VV/  **************************************************************)
(*    //   *    This file is distributed under the terms of the         *)
(*         *     GNU Lesser General Public License Version 2.1          *)
(*         *     (see LICENSE file for the text of the license)         *)
(************************************************************************)

Require Import Ltac2.Init.

Ltac2 Type t := constant.

Ltac2 @ external equal : constant -> constant -> bool := "rocq-runtime.plugins.ltac2" "constant_equal".
(** Constants obtained through module aliases or Include are not
    considered equal by this function. *)

Ltac2 @external print : t -> message
  := "rocq-runtime.plugins.ltac2" "constant_print".
(** Print the constant using the shortest qualified identifier which refers to it.
    Does not avoid variable names in the current or global environment. *)
